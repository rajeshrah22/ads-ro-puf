*run oscillator
.include ring_oscillator_0.cir
.include ring_oscillator_1.cir
.include ring_oscillator_2.cir
.include ring_oscillator_3.cir
.include ring_oscillator_4.cir
.include ring_oscillator_5.cir
.include ring_oscillator_6.cir
.include ring_oscillator_7.cir
.include nand.cir
.include inverter.sp

.global vdd
.global vss
VDD vdd 0 dc 1.2v
VSS vss 0 dc 0v

VEN en 0 pwl 0n 0v 4n 0v 5n 1v 100n 1v

.temp 13.5

XRO0 en out0 ring_oscillator_0
XRO1 en out1 ring_oscillator_1
XRO2 en out2 ring_oscillator_2
XRO3 en out3 ring_oscillator_3
XRO4 en out4 ring_oscillator_4
XRO5 en out5 ring_oscillator_5
XRO6 en out6 ring_oscillator_6
XRO7 en out7 ring_oscillator_7

.control
  set wr_vecnames
  set wr_singlescale

  alter VDD dc = 1.2
  set temp = 13.5
  tran 10p 100n
  run
  linearize
  wrdata all-1_2V-13_5C.csv all
  reset

  alter VDD dc = 1.2
  set temp = 27
  tran 10p 100n
  run
  linearize
  wrdata all-1_2V-27C.csv all
  reset

  alter VDD dc = 1.2
  set temp = 54
  tran 10p 100n
  run
  linearize
  wrdata all-1_2V-54C.csv all
  reset

  alter VDD dc = 1.5
  set temp = 27
  tran 10p 100n
  run
  linearize
  wrdata all-1_5V-27C.csv all
  reset

  alter VDD dc = 1.0
  set temp = 27
  tran 10p 100n
  run
  linearize
  wrdata all-1V-27C.csv all
  reset
.endc

*.control
*tran 10p 100n
*run
**save v(e) v(out0) v(out1) v(out2) v(out3) v(out4) v(out5) v(out6) v(out7)
*linearize
*set wr_vecnames
*set wr_singlescale
*wrdata all-1V_13_5C.csv all
**v(out7)
*.endc

.end
